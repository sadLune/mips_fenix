library IEEE;
use IEEE.STD_LOGIC_1164.all;

package blocks is
	type word_block is array (15 downto 0) of std_logic_vector(31 downto 0);
end package;
